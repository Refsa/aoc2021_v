module aoc11

pub struct AOC11 { }

pub fn (aoc AOC11) run_p1(input []string) ?u64 {
	return 0
}

pub fn (aoc AOC11) run_p2(input []string) ?u64 {
	return 0
}