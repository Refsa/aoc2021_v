module aoc8

pub struct AOC8 {}

pub fn (aoc AOC8) run_p1(input []string) ?u64 {
	return 0
}

pub fn (aoc AOC8) run_p2(input []string) ?u64 {
	return 0
}